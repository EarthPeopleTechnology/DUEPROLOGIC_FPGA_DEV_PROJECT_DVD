library verilog;
use verilog.vl_types.all;
entity i2c_slave_comms is
    generic(
        IDLE            : integer := 0;
        I2C_START       : integer := 1;
        READ_ADDRESS    : integer := 2;
        DECODE_RW       : integer := 3;
        CHECK_READ_WRITE: integer := 4;
        WRITE_BYTE      : integer := 5;
        WRITE_ACK       : integer := 6;
        WRITE_ACK_DELAY : integer := 7;
        READ_BYTE       : integer := 8;
        READ_ACK        : integer := 9;
        READ_ACK_DELAY  : integer := 10;
        I2C_STOP        : integer := 11;
        I2C_IDLE_STATE  : integer := 0;
        I2C_DATA_LOW_STATE: integer := 1;
        I2C_CLOCK_LOW_STATE: integer := 2;
        I2C_START_DETECT_STATE: integer := 3;
        I2C_ACK_DONE_STATE: integer := 4;
        I2C_CLOCK_HIGH_STATE: integer := 5;
        I2C_DATA_HIGH_STATE: integer := 6;
        I2C_WRITE_CLOCK_LOW_STATE: integer := 7;
        I2C_WRITE_DATA_LOW_STATE: integer := 8;
        I2C_STOP_DETECT_STATE: integer := 9;
        I2C_START_STOP_COUNT: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0);
        I2C_ERROR_COUNT : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1);
        I2C_WAIT_BYTE_COUNT: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1);
        DEVICE_ADDRESS  : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0)
    );
    port(
        CLK             : in     vl_logic;
        RESET           : in     vl_logic;
        IIC_DATA        : inout  vl_logic;
        IIC_CLOCK       : in     vl_logic;
        SERIAL_IIC_TRANSMIT_DATA_IN: in     vl_logic_vector(7 downto 0);
        SERIAL_IIC_TRANSMIT_ENA_OUT: out    vl_logic;
        SERIAL_IIC_TRANSMIT_RDY_IN: in     vl_logic;
        SERIAL_IIC_RECEIVE_DATA_OUT: out    vl_logic_vector(7 downto 0);
        SERIAL_IIC_RECEIVE_ENA_IN: in     vl_logic;
        SERIAL_IIC_RECEIVE_RDY_OUT: out    vl_logic;
        ERROR_OUT       : out    vl_logic_vector(7 downto 0);
        TEST_BUS_OUT    : out    vl_logic_vector(11 downto 0);
        STATE_OUT       : out    vl_logic_vector(3 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of IDLE : constant is 1;
    attribute mti_svvh_generic_type of I2C_START : constant is 1;
    attribute mti_svvh_generic_type of READ_ADDRESS : constant is 1;
    attribute mti_svvh_generic_type of DECODE_RW : constant is 1;
    attribute mti_svvh_generic_type of CHECK_READ_WRITE : constant is 1;
    attribute mti_svvh_generic_type of WRITE_BYTE : constant is 1;
    attribute mti_svvh_generic_type of WRITE_ACK : constant is 1;
    attribute mti_svvh_generic_type of WRITE_ACK_DELAY : constant is 1;
    attribute mti_svvh_generic_type of READ_BYTE : constant is 1;
    attribute mti_svvh_generic_type of READ_ACK : constant is 1;
    attribute mti_svvh_generic_type of READ_ACK_DELAY : constant is 1;
    attribute mti_svvh_generic_type of I2C_STOP : constant is 1;
    attribute mti_svvh_generic_type of I2C_IDLE_STATE : constant is 1;
    attribute mti_svvh_generic_type of I2C_DATA_LOW_STATE : constant is 1;
    attribute mti_svvh_generic_type of I2C_CLOCK_LOW_STATE : constant is 1;
    attribute mti_svvh_generic_type of I2C_START_DETECT_STATE : constant is 1;
    attribute mti_svvh_generic_type of I2C_ACK_DONE_STATE : constant is 1;
    attribute mti_svvh_generic_type of I2C_CLOCK_HIGH_STATE : constant is 1;
    attribute mti_svvh_generic_type of I2C_DATA_HIGH_STATE : constant is 1;
    attribute mti_svvh_generic_type of I2C_WRITE_CLOCK_LOW_STATE : constant is 1;
    attribute mti_svvh_generic_type of I2C_WRITE_DATA_LOW_STATE : constant is 1;
    attribute mti_svvh_generic_type of I2C_STOP_DETECT_STATE : constant is 1;
    attribute mti_svvh_generic_type of I2C_START_STOP_COUNT : constant is 1;
    attribute mti_svvh_generic_type of I2C_ERROR_COUNT : constant is 1;
    attribute mti_svvh_generic_type of I2C_WAIT_BYTE_COUNT : constant is 1;
    attribute mti_svvh_generic_type of DEVICE_ADDRESS : constant is 1;
end i2c_slave_comms;
