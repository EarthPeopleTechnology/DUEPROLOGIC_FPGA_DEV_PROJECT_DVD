library verilog;
use verilog.vl_types.all;
entity EPT_4CE6_AF_D1_Top is
    generic(
        GLOBAL_RESET_COUNT: vl_logic_vector(0 to 11) := (Hi1, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0);
        TRANSFER_HOST_IDLE: integer := 1;
        TRANSFER_HOST_LOOPBACK_START: integer := 2;
        TRANSFER_HOST_LOOPBACK_COMPLETE: integer := 3;
        BLOCK_COUNT_16  : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0);
        BLOCK_LOOPBACK_IDLE: integer := 1;
        BLOCK_LOOPBACK_INIT: integer := 2;
        FIFO_EN_HIGH    : integer := 3;
        FIFO_EN_LOW     : integer := 4;
        BLK_TRANSFER_OUT_IDLE: integer := 1;
        BLK_TRANSFER_OUT_COUNT: integer := 2;
        IDLE            : integer := 0;
        SELECT_MODE     : integer := 1;
        LOAD_REGISTER   : integer := 2;
        LOAD_LEDS       : integer := 3;
        WAIT_FOR_TIMER  : integer := 6;
        RANDOM_NUMBER   : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi1);
        SHIFT_LEFT      : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi1, Hi0);
        SHIFT_RIGHT     : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi1, Hi1);
        COUNT_UP        : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi0);
        COUNT_DOWN      : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi1);
        STATIC_VALUE    : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi0);
        TIMER_LOW_LIMIT : vl_logic_vector(0 to 23) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1)
    );
    port(
        aa              : in     vl_logic_vector(1 downto 0);
        bc_in           : in     vl_logic_vector(1 downto 0);
        bc_out          : out    vl_logic_vector(2 downto 0);
        bd_inout        : inout  vl_logic_vector(7 downto 0);
        XIO_1           : out    vl_logic_vector(7 downto 0);
        XIO_2           : out    vl_logic_vector(2 downto 0);
        XIO_2_IN        : in     vl_logic_vector(4 downto 0);
        XIO_3           : out    vl_logic_vector(7 downto 0);
        XIO_4           : out    vl_logic_vector(7 downto 0);
        XIO_5           : out    vl_logic_vector(7 downto 0);
        XIO_6           : out    vl_logic_vector(7 downto 0);
        XIO_7           : in     vl_logic_vector(5 downto 0);
        RESET           : out    vl_logic;
        UBA             : in     vl_logic;
        UBB             : in     vl_logic;
        SD_DATA         : in     vl_logic_vector(3 downto 0);
        SD_CMD          : out    vl_logic;
        SD_CLK          : out    vl_logic;
        ULG             : out    vl_logic;
        ULY             : out    vl_logic;
        ULO             : out    vl_logic;
        ULR             : out    vl_logic;
        LED             : out    vl_logic_vector(3 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of GLOBAL_RESET_COUNT : constant is 1;
    attribute mti_svvh_generic_type of TRANSFER_HOST_IDLE : constant is 1;
    attribute mti_svvh_generic_type of TRANSFER_HOST_LOOPBACK_START : constant is 1;
    attribute mti_svvh_generic_type of TRANSFER_HOST_LOOPBACK_COMPLETE : constant is 1;
    attribute mti_svvh_generic_type of BLOCK_COUNT_16 : constant is 1;
    attribute mti_svvh_generic_type of BLOCK_LOOPBACK_IDLE : constant is 1;
    attribute mti_svvh_generic_type of BLOCK_LOOPBACK_INIT : constant is 1;
    attribute mti_svvh_generic_type of FIFO_EN_HIGH : constant is 1;
    attribute mti_svvh_generic_type of FIFO_EN_LOW : constant is 1;
    attribute mti_svvh_generic_type of BLK_TRANSFER_OUT_IDLE : constant is 1;
    attribute mti_svvh_generic_type of BLK_TRANSFER_OUT_COUNT : constant is 1;
    attribute mti_svvh_generic_type of IDLE : constant is 1;
    attribute mti_svvh_generic_type of SELECT_MODE : constant is 1;
    attribute mti_svvh_generic_type of LOAD_REGISTER : constant is 1;
    attribute mti_svvh_generic_type of LOAD_LEDS : constant is 1;
    attribute mti_svvh_generic_type of WAIT_FOR_TIMER : constant is 1;
    attribute mti_svvh_generic_type of RANDOM_NUMBER : constant is 1;
    attribute mti_svvh_generic_type of SHIFT_LEFT : constant is 1;
    attribute mti_svvh_generic_type of SHIFT_RIGHT : constant is 1;
    attribute mti_svvh_generic_type of COUNT_UP : constant is 1;
    attribute mti_svvh_generic_type of COUNT_DOWN : constant is 1;
    attribute mti_svvh_generic_type of STATIC_VALUE : constant is 1;
    attribute mti_svvh_generic_type of TIMER_LOW_LIMIT : constant is 1;
end EPT_4CE6_AF_D1_Top;
